module alu32(sum,a,b,status,gin,stswrite);//ALU operation according to the ALU control line values
output [31:0] sum;
input [31:0] a,b; 
input [2:0] gin;//ALU control line
reg [31:0] sum;
reg [31:0] less;
output[2:0] status;
reg [2:0] status;
input stswrite;
always @(a or b or gin or stswrite)
begin
	case(gin)
	3'b010:
	begin
		sum=a+b; 		//ALU control line=010, ADD
		if(stswrite)
		begin
			status[0]=(sum[31] & ~a[31] & ~b[31]) | (~sum[31] & a[31] & b[31]); // overflow
		end
	end
	3'b110:
	begin
		sum=a+1+(~b);	//ALU control line=110, SUB
		if(stswrite)
		begin
			status[0]= (~sum[31]&a[31]&(~b[31]))|(sum[31]&~a[31]&b[31]); // overflow
		end
	end
	3'b111: begin less=a+1+(~b);	//ALU control line=111, set on less than
			if (less[31]) sum=1;	
			else sum=0;
		  end
	3'b000: sum=a & b;	//ALU control line=000, AND
	3'b001: sum=a|b;		//ALU control line=001, OR
	3'b101: sum=a<<b;
	default: sum=31'bx;	
	endcase
	
	if(stswrite)
	begin
		status[2]=~(|sum); // zero
		status[1]=sum[31]; // negative
		status[0]=(sum[31] & ~a[31] & ~b[31]) | (~sum[31] & a[31] & b[31]); // overflow
	end
end
endmodule
